BZh91AY&SY>F` G_�Ryg���w������`�      !&�ȍ &���40���L�1M00&�#��M C��4b�` `M0F	��� 0�2h�14�@��`�M4 a2dшbi���4�&&�h �I# LF��e2�4�C�=MO9�(�$���%�	&�s�I�O��]Y�c��S��������Ҙ��d�n���t����ukIb��R�%��K�&5!qI��&J)_�S�Q�\ԌJF���gm��>�g���V?�E��;��y�=�{߃Zض�4���
�3�b���(�K5�覟���i�i��e�Գ�cO9��a���p�{��%ZNg�t�_S�ly������k'�\v�6�9e�g��ϑ �z��qѷuU���)���}?G�Q���~1��~��EIJ��Q2�2:��t��ڋ�̮�{V&ơ�#3�Gf���G�P��P�R������U��ђ�Z�^�j��h[���X�R�b��;r��p�/��R�i�V���*���0V�-W���k��U1����]�=d����pX��V��������h�.��G��=3��=T��}#�����\�]ms��V%5�^�l�3*K�0�)1��5S�u��aQU�j�2�=��Ufmf��efQ��´�Uc�9�UUw���6lZM��Us�R��s̓��,Z� �]Ja	�������N�ο�}�0��[���F6����CFJm�4���r���UV~�GSͬ[����ס������m��?�9�?����c����bO懬e�G��H�EǶ~�<Ng�s��'V��b���<���u~S�6Z�.�6~�uƱNRO���>w�p]g��T��-{Bь��mSX�Ĩc�Lx��p�Y��H0Jg���)u�0�a��h�F���C�qFf�^R^��xV����)L���v�Tw��f,�8L/��E����͖Щb������M]qh���6����c;]{
��uG"�W�|�dx��a��⪊vY2{[�b�_]��ԆS�=���uCr�%�d*<c"y�u*R�<1��;�t�F����v��T�Bl�&�9���+;��N���u�;YO���q���k.�|�����Y�6I�r��S��c����oh�p��1�:
��9��|�>��
e��i;J��q�j�7g�j4=?f��4<S����d��YR�J)��T��K��#�X�6�眙��"�~��#3�ԗ����/RҬX�*vJKv��7��4V��}$�ţH�Z�Ō44�4iF;%썒L/����J�b�K����LC��R�w��0����i���opsk�)89NQywE�ENxti�v�����>ؓ���誴��s}�9�|Ws�.s�ުO��H�B��n��R,.P���<;�h�v���&ý�(k��r��H�;yֻ�1X�YE�a\�^3y���݋��y&�w�;Le�ʪ���gG�s'E�2�m0:�9�ݛ�a�W!��UͺYG�^-96�!Ý�_��I#f�.xP���E���1N��T�Z�}�[��拶��W�8�N��F�*I��,�*;['��������5J�?*C�s{z"7���ܑN$��� 