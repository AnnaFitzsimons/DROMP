BZh91AY&SY^�N �߀Ryg����������`|�ɠȹs� �+V� �#��  �@ �� 8���  0�2d�0��FLC �d �4ɓ�CA&��<hЦG��F�h�& �  �CIOe#�i��OP=A�4  4d�h(!2�cD�ѦB������d�����M4�pRFjC�0B��D�A:,���Y��٩��FA͝��#��X�>'/B[)�N���JN���#[��B�ix@��
�� �lE\�%у�R�]���%>��F�p�8F }YSl�/���'�ݯO~?�ͩ�Оg/�A�<mg<��0+o�+X3�Yrl��q� �Zҩe�cm'�u/Jke��MRj+���.7��j��R�J�(r.q25-��on}<�k����rMu�ց�G�8p
_�-M���r�|�`_"n7a|D����v�KӯpC�0�e�6E�y���6�"�V��pS��<�+�)�C��x�)u/��#p��,8��`�.[E��HC%�)�<�u�t� �Hs�&'�(9��h�-ƍLM�G0ֆ��o
J���Zб�3
��o��ln�(���OD�	�MDꄣ�mEM2��-*�����a�s^�7�u�5}Ii1h��	A�����ҷ�t�6U�/f��ThxQ��,��KU�Kʘ�����
a��4Ѩ�0񌒎.��Dɘ���əV�ن©iЅ�"�\� ��uUv��)|�$���H^gr� ��	B�AGn�����]bhC�K22������S_�qڼ(���P	�_4�h�[������A��/����fL9��\8����L�a�Ȱ���w�6��z��"w�� 0���V�� �㷧�mC��x�< Z� I�醷��d��G�^�&����Pnex��հ�5n�Ze&N�`{��}<����}�2����_��Z[1�B���D�m���!!�lJ'���c¢�I�66��Nz�z
{F���;��מÖ'xsS�0�Z�
�J�e=1�sr���v�W��=m<�!���Q�l0$R�Q�GJb(j��� F�L�	d��L2�(�:[<Y�I��I�h|���Ѡ�����sÑ$��.�`��;X�\�V��"V�M�c)�CPBt	Ԙ+�W6�a A����uB1/dV�:o� ����5o���h���'N$��n�s'8á��k9�C��{�|	�;<�s���K�Ɲ���Z��1j8�:9�<����D%��tA�pj�� Adk$�J�0�� ���� �>�~ce�b������8�)qQ�$`����#!`,D&��1����q Z����=W�8��2���Qj�؆	-j
�0d+KK}� ���-j��H$�HRl|���e�r2 �6�0&�o�����S��	�e+�.�Y�!�v�~���}�6�]����k�� ��;N&���QCs�8|,��ט�CX�G� {�=RP��N��6~��=��,�b��j<|���Y�T�� �`�&jQ�Y@j0�}}xc���h/Ϣ�3��i����"��f�*��80���H�sw܉�_/gML�Ҫ�'���FX�3HI]&[8?qկ_�����8Á�*�Xx+ۣ����GF�n�,tM��ء@�ϋ�������l�ݫ�z�?#��D}��e���y�>D�CF=e��ciҎ��<���
�����e�4ε
�Zƅ��c��!�u{���lp�ڌ`�1ߨ����H�
��)�