BZh91AY&SY��J %߀Ryg���g�����`	}�hP �)*� ��2dшbi���4�&&�h ��Hh     M4 8ɓF!���`��i�q�&�CL	��14�@D��S*{R?)6�OT�2~�~��OSdi�'��4�  )�Si�&چ�?Tb0ѣMN"�"0|3�`�74Dɴ������X(�;51�I��*��y���XA�I'	��K�P��CYS�p, ����7�����~�
�B�F�b�ɉ��J�X?�m'(�!���u�)�!���g����ߎ/�uli�=�Y��Al%!��I������<�ī�`��-$++Ķ��6�b
tR�#�e��6F�r�	j��Q W� .���8p���B�L)l�`X�Ά��3��Ӗ^������ϕ�˘|��|��ƯZZ��(�}~�Cn v'w	��x���ZrG���_�`B���y�N�o �u� �۰���ƞ���f�6�w�ӄr�wK@�\��8E0S��p _��<���I ɉ� ��@Т�\Y>����^��9d.�u�$MO>��q-ΚaX��������i�9K�HU���I0��X��fc�b��`���β���
?{$8�FJ�I$�I$��e6#I���O!<w�m��n�p��KC#N2��a �A��`av�24����?]c�!�	�@�/������B��cL���L���I$%9;ca3	�@͊���JOc�$l���@�R�l�I��ki��e��~��Nn����!��J��23@5�R*���<����ʛo�Ҩ"��1����Ԗw���(�#l9�&��RLL������=�Wv8;��hknuR����\p������^���A�-��'�! W>�	�]=j�Do/�0�� J��_��PP`t�pz��;����%��S�9�{ѻ:����������˴�@����M�I�߉@��g��"����2{-]@��!?��S�w�C8i���Mɖ�Z��zZ����4O���\��#''7��J=c}�]έ��[�!�B�Q�D('��egztﱎ�
88�4J5Y	pS�kXU�)���`ȥ!M4��� PX5.>��.�0ccc�,�>I���B��q�\C����2N`v'>�c������N�'H���H���^.&�U^~yJ{�1z�����ZۄB��;��x%��P���`��֗��l�HGƇ�c$�xp.�X�U��8S�>��>���S��F���{�y��q�纬h��ɚo��G6Ӹ�2�zfC�N��ۙ���FâV���F���C*�7q����_����7�&�v��G��G0� y���<��p h�?' rC�p�4@"OՑ�0b���
VݼC��	���n�����
u��"�&��
-N��� �� J

v�i�B����3�2m�))3%Ss��i��ffA�P���t�z��H�v���s�f�Ⱥ�����C���GqJ����0���9?.N���a��Q�~=�aOC�9�w
X����uk�>���#��@�#o?l�q�m�F����{O2�7F�wǧ�����3�J)��\��HŊ��b4����-ݙ��>� ��N
��b��䆣����"�ǣ��Gn��
�L:�8���s������>�MK��;��d̄�烌I�B�j��$����wc����3�z@�=���3��M0J�_�gW�e����u1kt�p-��(=��tn�; �49tp���#~~�����	���`R�~�0�k�ښ�Sߵ�ϼ�-�(�c����w��hv���٭�@��E�������HC-�m�����ь�9r���.�p�!�;x�